package Parameter_Definitions;

	parameter NBits = 8; //8

endpackage
