//import Parameter_Definitions::*;

module DIVISOR
(
	//Inputs			
	input clk,
	input rst,										
	input enable,
	input [15:0]Data,
	output [15:0]Result,
	output [15:0]Residue,//negated_shift_enable Tells you when it has finished so it stops the shifting
	output ready
	);


endmodule