package definitions; 

	parameter VERSION = "1.2";
	parameter NBits = 8;
endpackage	