package Parameter_Definitions;

	parameter NBits = 7;

endpackage
